LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY Bus_Arbiter IS

  -------------------------------------------------------------------------------
  --                             Port Declarations                             --
  -------------------------------------------------------------------------------
  PORT (
    -- Inputs
    clk               : IN STD_LOGIC;
    reset_n           : IN STD_LOGIC;
    cpu_0_address     : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
    cpu_0_bus_enable  : IN STD_LOGIC;
    cpu_0_byte_enable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    cpu_0_rw          : IN STD_LOGIC;
    cpu_0_write_data  : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    cpu_1_address     : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
    cpu_1_bus_enable  : IN STD_LOGIC;
    cpu_1_byte_enable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    cpu_1_rw          : IN STD_LOGIC;
    cpu_1_write_data  : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    -- Outputs
    cpu_0_acknowledge : OUT STD_LOGIC;
    cpu_0_read_data   : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    cpu_1_acknowledge : OUT STD_LOGIC;
    cpu_1_read_data   : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
  );
END Bus_Arbiter;

ARCHITECTURE Bus_Arbiter_rtl OF Bus_Arbiter IS

  --The Ram controller is taken from part 1. it is an interface from the bus bridge to the RAM

  COMPONENT RAM_controller IS
    PORT (
      clk     : IN STD_LOGIC := 'X'; -- clk
      reset_n : IN STD_LOGIC := 'X'; -- reset_n
      ---- Bridge Interface 
      bridge_acknowledge : OUT STD_LOGIC := 'X';                                 -- acknowledge
      bridge_irq         : OUT STD_LOGIC := 'X';                                 -- irq
      bridge_address     : IN STD_LOGIC_VECTOR(10 DOWNTO 0);                     -- address
      bridge_bus_enable  : IN STD_LOGIC;                                         -- bus_enable
      bridge_byte_enable : IN STD_LOGIC_VECTOR(1 DOWNTO 0);                      -- byte_enable
      bridge_rw          : IN STD_LOGIC;                                         -- rw (0 = write, 1= read)
      bridge_write_data  : IN STD_LOGIC_VECTOR(15 DOWNTO 0);                     -- write_data
      bridge_read_data   : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => 'X'); -- read_data
      ---- RAM interface
      ram_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      ram_data    : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      ram_wren    : OUT STD_LOGIC;
      ram_q       : IN STD_LOGIC_VECTOR (15 DOWNTO 0));
  END COMPONENT;

  --the external RAM is generated by Altera MegaWizard Plug-in Manager	
  COMPONENT external_RAM IS
    PORT (
      address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
      clock   : IN STD_LOGIC := '1';
      data    : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      wren    : IN STD_LOGIC;
      q       : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
  END COMPONENT;

  --the arbiter is a state machine so define the states here
  TYPE state_type IS (IDLE, CPU_0, CPU_1);
  SIGNAL current_state, next_state : state_type;

  -------------------------------------------------------------------------------
  --                 Internal Wires                                            --
  -------------------------------------------------------------------------------
  -- Internal Wires

  SIGNAL bus_enable_both             : STD_LOGIC_VECTOR(1 DOWNTO 0);
  SIGNAL acknowledge, bus_enable, rw : STD_LOGIC;
  SIGNAL read_data, write_data       : STD_LOGIC_VECTOR(15 DOWNTO 0);
  SIGNAL address                     : STD_LOGIC_VECTOR(10 DOWNTO 0);
  SIGNAL byte_enable                 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  SIGNAL irq                         : STD_LOGIC;

  SIGNAL ram_address_int : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL ram_data_int    : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL ram_wren_int    : STD_LOGIC;
  SIGNAL ram_q_int       : STD_LOGIC_VECTOR (15 DOWNTO 0);

BEGIN

  -- create a signal to indicate which bridge has been enabled
  bus_enable_both <= cpu_0_bus_enable & cpu_1_bus_enable;

  -------------------------------------------------------------------------------
  --                         Finite State Machine                              --
  -------------------------------------------------------------------------------
  sync : PROCESS (clk, reset_n)
  BEGIN
    IF (reset_n = '0') THEN
      current_state <= IDLE;
    ELSIF (clk'event AND clk = '1') THEN
      current_state <= next_state;
    END IF;
  END PROCESS;
  -------------------------------------------------------------------------------
  --                            Combinational Logic                            --
  -------------------------------------------------------------------------------
  comb : PROCESS (current_state, bus_enable_both, bus_enable)
  BEGIN
    CASE(current_state) IS
      WHEN idle =>
      CASE (bus_enable_both) IS
        WHEN "10" =>
          next_state <= CPU_0;
        WHEN "01" =>
          next_state <= CPU_1;
        WHEN "11" =>
          --Need to arbitrate here
          --Determine an arbitration scheme so that the two processors are fairly
          --       given access to the bus
          next_state <= CPU_0;
        WHEN OTHERS =>
          next_state <= IDLE;
      END CASE;
      WHEN CPU_0 =>
      IF (bus_enable = '0') THEN
        next_state <= IDLE;
      ELSE
        next_state <= CPU_0;
      END IF;
      WHEN CPU_1 =>
      IF (bus_enable = '0') THEN
        next_state <= IDLE;
      ELSE
        next_state <= CPU_1;
      END IF;
      WHEN OTHERS =>
      next_state <= IDLE;
    END CASE;
  END PROCESS;
  --this process assigns all of the signals based on which bridge is selected
  --Note - it is not the best coding style to use one process for all the 
  --  outputs (j. christman)

  PROCESS (current_state, cpu_0_bus_enable, cpu_0_byte_enable, cpu_0_rw,
    cpu_0_address, cpu_0_write_data, cpu_1_bus_enable, cpu_1_byte_enable, cpu_1_rw,
    cpu_1_address, cpu_1_write_data) IS
  BEGIN
    CASE (current_state) IS
      WHEN CPU_0 =>
        bus_enable        <= cpu_0_bus_enable;
        byte_enable       <= cpu_0_byte_enable;
        rw                <= cpu_0_rw;
        address           <= cpu_0_address;
        write_data        <= cpu_0_write_data;
        cpu_0_acknowledge <= acknowledge;
        cpu_0_read_data   <= read_data;
        cpu_1_acknowledge <= '0';
        cpu_1_read_data   <= (OTHERS => '0');

      WHEN OTHERS =>
        bus_enable        <= cpu_1_bus_enable;
        byte_enable       <= cpu_1_byte_enable;
        rw                <= cpu_1_rw;
        address           <= cpu_1_address;
        write_data        <= cpu_1_write_data;
        cpu_0_acknowledge <= '0';
        cpu_0_read_data   <= (OTHERS => '0');
        cpu_1_acknowledge <= acknowledge;
        cpu_1_read_data   <= read_data;

    END CASE;
  END PROCESS;
  -------------------------------------------------------------------------------
  --                              Internal Modules                             --
  -------------------------------------------------------------------------------
  u1 : RAM_controller
  PORT MAP
  (
    clk     => clk,
    reset_n => reset_n,
    ---- Bridge Interface 
    bridge_acknowledge => acknowledge,
    bridge_irq         => irq,
    bridge_address     => address,
    bridge_bus_enable  => bus_enable,
    bridge_byte_enable => byte_enable,
    bridge_rw          => rw,
    bridge_write_data  => write_data,
    bridge_read_data   => read_data,
    ---- RAM interface
    ram_address => ram_address_int,
    ram_data    => ram_data_int,
    ram_wren    => ram_wren_int,
    ram_q       => ram_q_int
  );

  u2 : external_RAM
  PORT MAP
  (
    address => ram_address_int,
    clock   => clk,
    data    => ram_data_int,
    wren    => ram_wren_int,
    q       => ram_q_int
  );

END Bus_Arbiter_rtl;
