LIBRARY ieee; 
USE ieee.std_logic_1164.all; 
USE ieee.numeric_std.all;
USE ieee.std_logic_unsigned.all; 

LIBRARY WORK;
USE WORK.servo_controller_pkg.ALL;

ENTITY top IS
PORT ( 	
  CLOCK_50  : IN STD_LOGIC; 					-- 50MHz clock
  reset     : IN STD_LOGIC;
  write    : IN  STD_LOGIC;
  SW 	    : IN STD_LOGIC_VECTOR(9 DOWNTO 0);	-- Switch inputs
  writedata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
  address   : IN STD_LOGIC;
  LEDR	    : OUT STD_LOGIC_VECTOR(9 DOWNTO 0); -- LED outputs
  irq       : OUT STD_LOGIC;					-- IRQ output
  outwave   : OUT STD_LOGIC
  ); 
END top; 

ARCHITECTURE Structure OF top IS

  SIGNAL reset_n  : STD_LOGIC := '0';
  
  SIGNAL key0_d1  : STD_LOGIC;
  SIGNAL key0_d2  : STD_LOGIC;
  SIGNAL key0_d3  : STD_LOGIC;
  
  SIGNAL max_angle : UNSIGNED(31 DOWNTO 0);
  SIGNAL min_angle : UNSIGNED(31 DOWNTO 0);
  
BEGIN
-- Instantiate the Nios II system entity generated by the SOPC Builder 

  ----- Synchronize Keys
  synchReset_proc : PROCESS (CLOCK_50)
  BEGIN
    IF (RISING_EDGE(CLOCK_50)) THEN
	  key0_d1 <= reset;
      key0_d2 <= key0_d1;
      key0_d3 <= key0_d2;
    END IF;
  END PROCESS synchReset_proc;

  reset_n 	  <= key0_d3;
  
  servo_top : servo_controller
  GENERIC MAP (
    max_angle => to_unsigned(1000000, 32),
    min_angle => to_unsigned(50000, 32)
	)
  PORT MAP(
    CLOCK_50 => CLOCK_50,
    reset => reset_n,
    write => write,
    writedata => writedata,
	address => address,
    irq => irq,
    LEDR => LEDR,
	outwave => outwave
    );

END Structure;
