
module nios_system (
	clk_clk,
	reset_reset_n,
	servo_controller_ext_out_wave);	

	input		clk_clk;
	input		reset_reset_n;
	output		servo_controller_ext_out_wave;
endmodule
